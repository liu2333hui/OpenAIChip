`define	REQUIRED_PES	16
`define	MAX_WEI_PRECISION	16
`define	MAX_ACT_PRECISION	16
`define	MIN_WEI_PRECISION	16
`define	MIN_ACT_PRECISION	16
`define	MAX_OUT_PRECISION	16
`define	MIN_OUT_PRECISION	0
`define	MAX_ELEMENT_UNITS	0
`define	MAX_WEI_PRECISION_INT	16
`define	MIN_WEI_PRECISION_INT	16
`define	MAX_ACT_PRECISION_INT	16
`define	MIN_ACT_PRECISION_INT	16
`define	MAX_OUT_PRECISION_INT	16
`define	MIN_OUT_PRECISION_INT	16
`define	MAX_WEI_PRECISION_FP	0
`define	MIN_WEI_PRECISION_FP	0
`define	MAX_ACT_PRECISION_FP	0
`define	MIN_ACT_PRECISION_FP	0
`define	MAX_PRECISION_FP	0
`define	MAX_PSUM_PRECISION	32
`define	MAX_PSUM_PRECISION_INT	32
`define	MAX_PSUM_PRECISION_FP	0
`define	MAX_ACC_PRECISION	41
`define	MAX_ACC_PRECISION_INT	41
`define	MAX_ACC_PRECISION_FP	0
`define	CONV2D_OP	0
`define	LINEAR_OP	1
`define	TRANSFORMER_OP	2
`define	MAX_STRIDE	2
`define	MAX_KX	3
`define	MAX_KY	3
`define	MAX_X	128
`define	MAX_Y	128
`define	MAX_N	64
`define	MAX_I	64
`define	MAX_B	1
`define	MAX_PADDING_X	1
`define	MAX_PADDING_Y	1
`define	MAX_STRIDE_LOG	2
`define	MAX_KX_LOG	3
`define	MAX_KY_LOG	3
`define	MAX_X_LOG	8
`define	MAX_Y_LOG	8
`define	MAX_N_LOG	7
`define	MAX_I_LOG	7
`define	MAX_B_LOG	1
`define	MAX_PADDING_X_LOG	1
`define	MAX_PADDING_Y_LOG	1
`define	WEI_BUF_DATA	256
`define	ACT_BUF_DATA	64
`define	PSUM_BUF_DATA	192
`define	WEI_BUF_ROWS	8192
`define	WEI_BUF_ROWS_LOG2	13
`define	PSUM_BUF_ROWS	1024
`define	PSUM_BUF_ROWS_LOG2	10
`define	ACT_BUF_ROWS	16384
`define	ACT_BUF_ROWS_LOG2	14
`define	L2_WEI_BUF_ROWS	8192
`define	L2_WEI_BUF_ROWS_LOG2	13
`define	L2_ACT_BUF_ROWS	32768
`define	L2_ACT_BUF_ROWS_LOG2	15
