`define MAX_PRECISION 8
`define CLK_PERIOD 10
